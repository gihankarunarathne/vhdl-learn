----------------------------------------------------------------------------------
-- Company: UOM
-- Engineer: Gihan Karunarathne
-- 
-- Create Date:    13:03:09 08/21/2013 
-- Design Name: 
-- Module Name:    Priority_encoder - Behavioral 
-- Project Name:   tutorial I
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Priority_encoder is
end Priority_encoder;

architecture Behavioral of Priority_encoder is

begin

	

end Behavioral;

